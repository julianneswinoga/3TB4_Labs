module decoder (
	input [7:2] instruction,
	output br, brz, addi, subi, sr0, srh0, clr, mov, mova, movr, movrhs, pause
	);

assign br = (instruction[7:5] == 3'b100);
assign clr = (instruction[7:2] == 6'b011000);

//assign brz = (...);
//assign addi = (...);
//assign subi = (...);
//assign sr0 = (...);
//assign srh0 = (...);
//assign mov = (...);
//assign mova = (...);
//assign movr = (...);
//assign movrhs = (...);
//assign pause = (...);

endmodule
